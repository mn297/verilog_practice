module hello;
  initial 
    begin
      $display("Hello, WORLD!!!!");
      $finish ;
    end
endmodule